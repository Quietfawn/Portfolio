package uart_pkg;
  parameter int unsigned CLK_HZ = 100_000_000;
  parameter int unsigned BAUD   = 115200;
endpackage
